// python script nnet_verilog.py
// INPUT: filename.nnet
// OUTPUT: parsed filename.sv

/*
    Example:
    INPUT: filename.nnet


    OUTPUT: filename.sv
    -1.00006	e+00
    -1.00053	e+00
    -1.00315	e+00
    -1.00441	e+00
    ...
*?
